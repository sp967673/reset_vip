
`ifndef RESET_VIP_PKG
`define RESET_VIP_PKG

package reset_vip_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "reset_transaction.sv"
  `include "reset_driver.sv"
  `include "reset_monitor.sv"
  `include "reset_sequencer.sv"
  `include "reset_agent.sv"
  `include "reset_sequences.sv"

endpackage

`endif //RESET_VIP_PKG_SV
